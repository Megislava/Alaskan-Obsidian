module logicalOr(input a, b, output y);
	assign y = (a | b);
endmodule
